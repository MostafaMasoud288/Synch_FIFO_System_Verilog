package shared_pck;
integer error_count=0;
integer correct_count=0;
logic test_finished;
endpackage
